// Part 2 skeleton

module part2
	(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
        KEY,
        SW,
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0]
	);

	input			CLOCK_50;				//	50 MHz
	input   [9:0]   SW;
	input   [3:0]   KEY;

	// Declare your inputs and outputs here
	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	
	wire resetn;
	assign resetn = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.
	wire [2:0] colour;
	wire [7:0] x;
	wire [6:0] y;
	wire writeEn;

	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(colour),
			.x(x),
			.y(y),
			.plot(writeEn),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "black.mif";
			
	// Put your code here. Your code should produce signals x,y,colour and writeEn/plot
	// for the VGA controller, in addition to any other functionality your design may require.
    
    // Instansiate datapath
	// datapath d0(...);
	

    // Instansiate FSM control
    // control c0(...);
	combination c0(
		.clock(CLOCK_50),
		.resetn(resetn),
		.go(~KEY[3]),
		.display(~KEY[1]),
		.position_in(SW[6:0]),
		.color_in(SW[9:7]),
		.position_x(x),
		.position_y(y),
		.color_out(colour),
		.plot(writeEn)
		);
	 
	 
	 
endmodule

module datapath(
	input [6:0] position_in,
	input [2:0] color_in,
	input clk,
	input resetn,
	input ld_x, ld_y, draw,
	input [1:0] alu_x_op, alu_y_op,
	
	output reg [7:0] x_out,
	output reg [6:0] y_out,
	output reg [2:0] color_out
	);
	
	
	// input registers
	reg [7:0] x;
	reg [6:0] y;
	
	// output of the alu_x and alu_y
	reg [7:0] alu_x_out;
	reg [6:0] alu_y_out;
	
	
	// register x, y with respective logic
	always @(posedge clk) begin
		if (!resetn) begin
			x <= 8'b00000000;
			y <= 7'b0000000;
		end
		else begin
			if (ld_x) 
				x <= {1'b0, position_in};  //load alu_x_out if ld_alu_out is high, else load from position_in (user input)
			if (ld_y)
				y <= position_in;
		 end
	end
	
	// output result register
	always @(*) begin
		if (!resetn) begin
			x_out <= 8'b0;
			y_out <= 7'b0;
		end
		else begin 
			if (draw) begin
				x_out <= alu_x_out;
				y_out <= alu_y_out;
				color_out <= color_in;
			end
		end
	end

	
	// The ALU, we have two ALU, alu_x and alu_y
	always @(*)
	begin: ALU
		case (alu_x_op)
			default: alu_x_out <= {x[7:2], x[1:0] + alu_x_op};
		endcase
		
		case (alu_y_op)
			default: alu_y_out <= {y[6:2], y[1:0] + alu_y_op};
		endcase
	end
	
endmodule


module control(
	input clock,
	input resetn,
	input go, // load x and y
	input display, //draw the pixels
	
	output reg [1:0] alu_x_op,
	output reg [1:0] alu_y_op,
	output reg ld_x, ld_y, draw,
	output reg plot
	);
	
	reg [3:0] counter;
	reg [2:0] current_state, next_state;
	
	localparam  S_LOAD_X = 3'd0,
					S_LOAD_X_WAIT= 3'd1,
					S_LOAD_Y = 3'd2,
					S_LOAD_Y_WAIT = 3'd3,
					S_DISPLAY = 3'd4;
	
	
	
	always @(*)
	begin: states
		case (current_state)
			S_LOAD_X: next_state = go ? S_LOAD_X_WAIT : S_LOAD_X;
			S_LOAD_X_WAIT: next_state = go ? S_LOAD_X_WAIT : S_LOAD_Y;    // load x to register x
			S_LOAD_Y: next_state = go ? S_LOAD_Y_WAIT : S_LOAD_Y;
			S_LOAD_Y_WAIT: next_state = display ? S_DISPLAY  : S_LOAD_Y_WAIT;  // load y to register y
			S_DISPLAY: begin
				if (counter == 4'b1111) 
					next_state = S_LOAD_X;
				else 
					next_state = S_DISPLAY;
			end
			default: next_state = S_LOAD_X;
		endcase  // state table
	end

	
	
	// current state registers
	always @(posedge clock)
		 begin: state_FFs
			  if(!resetn)
					current_state <= S_LOAD_X;
			  else
					current_state <= next_state;
		 end // state_FFS
		 
	// Output logic aka all of our datapath control signals
	always @(*)
	begin: enable_signals
		// By default make all our signals 0
		ld_x = 1'b0;
		ld_y = 1'b0;
		alu_x_op = 2'b00;
		alu_y_op = 2'b00;
		draw = 1'b0;
		plot = 1'b0;
		
		case (current_state) 
			S_LOAD_X: begin
				ld_x <= 1'b1;
				end
			S_LOAD_Y: begin
				ld_y <= 1'b1;
				end
			S_DISPLAY: begin 
				ld_x <= 1'b1;
				ld_y <= 1'b1;
				alu_x_op <= counter[3:2];
				alu_y_op <= counter[1:0];
				draw <= 1'b1;
				plot <= 1'b1;
				end
			
		endcase
	end
	
	always @(posedge clock)
		if (!resetn) begin
			counter <= 4'b0000;
		end
		else if (current_state == 3'd4)
			begin
				if(counter == 4'b1111) begin
					counter <= 4'b0000;
					next_state <= S_LOAD_X;
				end
				else
					counter <= counter + 1'b1;
			end
	

endmodule

module combination(
	input clock,
	input resetn,
	input go,
	input display,
	input [6:0] position_in,
	input [2:0] color_in,
	 
	output [7:0] position_x,
	output [6:0] position_y,
	output [2:0] color_out,
	output plot
	);
	
	wire ld_x;
	wire ld_y;
	wire draw;
	wire [1:0] alu_x_op;
	wire [1:0] alu_y_op;

	
	datapath d0(
		.position_in(position_in),
		.color_in(color_in),
		.clk(clock),
		.resetn(resetn),
		.ld_x(ld_x),
		.ld_y(ld_y),
		.draw(draw),
		.alu_x_op(alu_x_op),
		.alu_y_op(alu_y_op),
		.x_out(position_x),
		.y_out(position_y),
		.color_out(color_out)
		);
	
	control c0(
		.clock(clock),
		.resetn(resetn),
		.go(go),
		.display(display),
		.draw(draw),
		.alu_x_op(alu_x_op),
		.alu_y_op(alu_y_op),
		.ld_x(ld_x),
		.ld_y(ld_y),
		.plot(plot)
		);
		
endmodule
		

	
	
	
